module adder_testbench;
    reg clk, rst, go;
    reg [3:0] A, B, C, D;
    wire [15:0] o_sum;

    adder

endmodule