module datapath (
    input clk,
    input rst,
    input [3:0] A, B, C, D,
    output reg [15:0] sum
);
    
endmodule