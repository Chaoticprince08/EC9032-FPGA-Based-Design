module controller (
    input clk,rst,
);
    
endmodule